`ifndef demux16
 `define demux16_v

`timescale 1ns/1ps

///////////////////////////////////////////////////////////////////////////////
//
// 16-BIT DEMULTIPLEXER WITH ENABLE
//
///////////////////////////////////////////////////////////////////////////////


module demux16(a, en, y);
   input [3:0] a;
	input en;
   reg [15:0]  y0;
   output [15:0] y;
   
   always @ (a) begin
      case (a)
	0: y0 = 16'b1111111111111110;
	1: y0 = 16'b1111111111111101;
	2: y0 = 16'b1111111111111011;
	3: y0 = 16'b1111111111110111;
	4: y0 = 16'b1111111111101111;
	5: y0 = 16'b1111111111011111;
	6: y0 = 16'b1111111110111111;
	7: y0 = 16'b1111111101111111;
	8: y0 = 16'b1111111011111111;
	9: y0 = 16'b1111110111111111;
	10: y0 = 16'b1111101111111111;
	11: y0 = 16'b1111011111111111;
	12: y0 = 16'b1110111111111111;
	13: y0 = 16'b1101111111111111;
	14: y0 = 16'b1011111111111111;
	15: y0 = 16'b0111111111111111;
      endcase // case (a)
   end // always @ (a)

   assign y = en == 1'b1 ? y0 : 16'b1111111111111111;
endmodule // demux16

`endif //  `ifndef demux16

// End of file.

