-------------------------------------------------------------------------------
--  File name: vcc.vhd
-------------------------------------------------------------------------------
--  Copyright (C) 1996, 1997  Free Model Foundry; http://www.FreeModelFoundry.com
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License version 2 as
--  published by the Free Software Foundation.
--
--  MODIFICATION HISTORY:
--
--  version: |  author:  | mod date: | changes made:
--    V1.0     R. Steele   97 APR 21   Initial release
--    V1.1     R. Steele   97 JUN 25   Added use vital
--------------------------------------------------------------------------------
--   PART DESCRIPTION:
-- 
--   Library:       SOURCES
--   Technology:    N/A
--   Part:          VCC
-- 
--   Description: Source of simulation value VCC -> std_logic '1'
-- 
--------------------------------------------------------------------------------
LIBRARY IEEE;   USE IEEE.std_logic_1164.ALL;
                USE IEEE.VITAL_primitives.all;
                USE IEEE.VITAL_timing.all;

--------------------------------------------------------------------------------
-- ENTITY DECLARATION
--------------------------------------------------------------------------------
ENTITY vcc IS
    port (    
            PWR   : OUT   std_logic := '1'  
         );

    ATTRIBUTE VITAL_level0 OF vcc : ENTITY IS TRUE;
END vcc;

--------------------------------------------------------------------------------
-- ARCHITECTURE DECLARATION
--------------------------------------------------------------------------------
ARCHITECTURE vhdl_behavioral OF vcc IS
    ATTRIBUTE VITAL_level1 OF vhdl_behavioral : ARCHITECTURE IS FALSE;
BEGIN
    PWR <= '1';

END vhdl_behavioral;
