///////////////////////////////////////////////////////////////////////////////
//
// THE DATA BUS INTERFACE (INCLUDING WAIT STATES)
//
// REDESIGNED IN 2019
//
// NOTES:
//
///////////////////////////////////////////////////////////////////////////////


`ifndef databus_v
`define databus_v

`include "buffer.v"
`include "flipflop.v"

`timescale 1ns/1ps

module databus (nreset, nhalt, clk3, clk4, t34,
		nmem, nio, nr, nwen,
		nws, nwaiting,
		ibus,
		nw, db);

   input 	nreset;
   input 	nhalt;
   input 	clk3;
   input 	clk4;
   input 	t34;
   input 	nmem;
   input 	nio;
   input 	nr;
   input 	nwen;
   inout 	nws;
   output 	nwaiting;

   inout [15:0] ibus;		// input & output!

   output 	nw;

   inout [15:0] db;		// input & output!

   wire 	nreset;
   wire 	nhalt;
   wire 	clk3;
   wire 	t34;
   wire 	nmem;
   wire 	nio;
   wire 	nr;
   wire 	nwen;
   tri1 	nws;		// Pulled up (may not be needed if Bus Hold is used)

   wire [15:0] 	ibus;
   
   wire 	nw;

   wire [15:0] 	db;

   // Wait states

   wire 	halt, nw0, nwaiting, nws_in_t34, nbusen;

   // The delays here are purposefully different, and all are much higher than
   // the maximum propagation delays for LVC family little gates.

   // nws_in_t34 ensures wait states are only requested during the last 50% of
   // the clock cycle.
   assign #7 nws_in_t34 = nws | t34;          // 74LVC1G32

   // Assign nWSTB to either CLK4 (original and tested configuration,
   // but with potential problems) or a custom, delayed
   // signal. (generated by a PLL clock doubler in hardware).
   reg 		clk4x8;
   // Generate a frequency 8× that of clk4 (using a PLL).
   always @ (negedge clk4) begin
      clk4x8 = 0;		// 0
      #31.25 clk4x8 = 1;

      #31.25 clk4x8 = 0;	// 1
      #31.25 clk4x8 = 1;

      #31.25 clk4x8 = 0;	// 2
      #31.25 clk4x8 = 1;

      #31.25 clk4x8 = 0;	// 3
      #31.25 clk4x8 = 1;
   end // always @ (negedge clk4)

   // Choose one assignment (JP3 on the BUS board).
   wire nwstb;
   //assign nwstb = clk4;
   assign #4 nwstb = clk4 | clk4x8;

   // The nW driver. The Microcode Sequencer can tri-state all its outputs when
   // nHALT is asserted, but we generate nW here, so we need to be able to tri-state it.
   assign #6 halt = ~nhalt;		      // 74LVC1G04
   //assign #8 nw0 = nwen | (wstb & nwaiting); // 74LVC1G0832
   // assign #8 nw0 = nwaiting & (nwen | clk4);
   assign #8 nw0 = nwaiting_delayed & (nwen | nwstb);
   assign #6 nw = halt ? 1'bz : nw0;	      // 74LVC1G125

   // The Wait State FF itself
   flipflop_74h #2.5 ff_ws (.nset(nws_in_t34), .d(1'b0), .clk(clk3), .nrst(nreset), .nq(nwaiting));

   // nwaiting must be deasserted after nwstb, but the rising edge of
   // nwstb can lead nwaiting's depending on jitter. If this condition
   // isn't satisfied, W# may glitch during wait states.
   wire nwaiting_delayed0, nwaiting_delayed;
   assign #4 nwaiting_delayed0 = nwaiting & nwaiting;
   assign #4 nwaiting_delayed = nwaiting & nwaiting_delayed0;

   assign #7 nbusen = nwaiting & nio & nmem; // 74LVC1G11

   // Connect the buses.
   buffer_245 buf_dblo (.a(ibus[7:0]),  .b(db[7:0]),  .dir(nr), .nen(nbusen));
   buffer_245 buf_dbhi (.a(ibus[15:8]), .b(db[15:8]), .dir(nr), .nen(nbusen));
   
endmodule // databus

`endif //  `ifndef databus_v

// End of file
